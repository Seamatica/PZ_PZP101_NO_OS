
module udp(
    input                rst_n       , //��λ�źţ��͵�ƽ��Ч
    
    input   wire [47:0]  board_mac,
    input   wire [31:0]  board_ip,
    input   wire [47:0]  des_mac,
    input   wire [31:0]  des_ip,
    input   wire [15:0]  board_port,
    input   wire [15:0]  des_port,    
    
    input                gmii_rx_clk , //KSZ9031_GMII��������ʱ��
    input                gmii_rx_en  , //KSZ9031_GMII����������Ч�ź�
    input        [7:0]   gmii_rxd    , //KSZ9031_GMII��������
    input                gmii_tx_clk , //KSZ9031_GMII��������ʱ��    
    output               gmii_tx_en  , //KSZ9031_GMII���������Ч�ź�
    output       [7:0]   gmii_txd    , //KSZ9031_GMII������� 
    output               rec_pkt_done, //��̫���������ݽ�������ź�
    output               rec_en      , //��̫�����յ�����ʹ���ź�
    output       [31:0]  rec_data    , //��̫�����յ�����
    output       [15:0]  rec_byte_num, //��̫�����յ���Ч�ֽ���    
    input                tx_start_en , //��̫����ʼ�����ź�
    input        [31:0]  tx_data     , //��̫������������  
    input        [15:0]  tx_byte_num , //��̫�����͵���Ч�ֽ���    
    output               tx_done     , //��̫����������ź�
    output               tx_req        //�����������ź�    
    );

//parameter  BOARD_MAC = 48'h00_00_99_00_33_11;     
//parameter  BOARD_IP  = {8'd192,8'd168,8'd1,8'd10};  
//parameter  DES_MAC   = 48'hff_ff_ff_ff_ff_ff;       
//parameter  DES_IP    = {8'd192,8'd168,8'd1,8'd11};

//wire define
wire          crc_en  ; //CRC��ʼУ��ʹ��
wire          crc_clr ; //CRC���ݸ�λ�ź� 
wire  [7:0]   crc_d8  ; //�����У��8λ����

wire  [31:0]  crc_data; //CRCУ������
wire  [31:0]  crc_next; //CRC�´�У���������

///////////////////////main code////////////////////////////////

assign  crc_d8 = gmii_txd;

//��̫������ģ��    
udp_rx u_udp_rx(
    .clk             (gmii_rx_clk ),        
    .rst_n           (rst_n       ),             
    .gmii_rx_en      (gmii_rx_en  ),                                 
    .gmii_rxd        (gmii_rxd    ),       
    .rec_pkt_done    (rec_pkt_done),      
    .rec_en          (rec_en      ),            
    .rec_data        (rec_data    ),          
    .rec_byte_num    (rec_byte_num),
    
    .board_mac       (board_mac),         //��������
    .board_ip        (board_ip )       
    );                                    

//��̫������ģ��
udp_tx u_udp_tx(
    .clk             (gmii_tx_clk),        
    .rst_n           (rst_n      ),             
    .tx_start_en     (tx_start_en),                   
    .tx_data         (tx_data    ),           
    .tx_byte_num     (tx_byte_num),    
    .crc_data        (crc_data   ),          
    .crc_next        (crc_next[31:24]),
    .tx_done         (tx_done    ),           
    .tx_req          (tx_req     ),            
    .gmii_tx_en      (gmii_tx_en ),         
    .gmii_txd        (gmii_txd   ),       
    .crc_en          (crc_en     ),            
    .crc_clr         (crc_clr    ),
    
    .board_mac       (board_mac),         //��������
    .board_ip        (board_ip ),
    .des_mac         (des_mac  ),
    .des_ip          (des_ip   ),
    .board_port      (board_port),
    .des_port        (des_port)            
    );                                      

//��̫������CRCУ��ģ��
crc32_d8   u_crc32_d8(
    .clk             (gmii_tx_clk),                      
    .rst_n           (rst_n      ),                          
    .data            (crc_d8     ),            
    .crc_en          (crc_en     ),                          
    .crc_clr         (crc_clr    ),                         
    .crc_data        (crc_data   ),                        
    .crc_next        (crc_next   )                         
    );

endmodule